// module av_cache_2w_v (Resetn, MEM_address, MEM_in, WR, Clock, MEM_out, Done);
module av_cache_2w_slave0_v (Resetn, MEM_address, MEM_in, WR, c0, c1,c2, MEM_out, Done);

// The address structure is: TAG=9-bit | Group=2-bit | Word=3-bit

parameter ma_max =    14,  // memory address width
          md_max =    14,  // memory data width 
		  ca_max =    6,   // cache address width {replace-bit, group-bits,word address bits} = 1+2+3=6
		  t_cnt_max = 3;   // words per block = 8 (=2^(3)) i.e. 3 bits. will be used to capture transfer count of words within a block
		  
parameter cam_addrs_max = 2, // | Group=2-bit| CAM address width, we have 4 locations so need only 2-bits to address them. 
          cam_arg_max =   9, // TAG=9-bit | CAM data width  = TAG size = 9-bits
		  cam_depth_max = 4; // total locations in CAM = number of groups (2^(2) = 4)

// Declare top module input and output ports //
input Resetn;  //Clock
input c0, c1, c2;
input WR;
input [ma_max-3:0] MEM_address;                    /* this is the address we receive from the CPU. 14-bit address, 
                                                      but we will only use 12-bit address to speedup the simulation. */
													  
/* MEM_address (memory address) = TAG=7-bit [11:5]| Group=2-bit [4:3]| Word=3-bit [2:0] */

input [md_max-1:0] MEM_in; // this the 14-bit data input

output [md_max-1:0] MEM_out; // this is the 14-bit data output 

output reg Done;
/*Means READ or WRITE ACCESS is complete, i.e. the output is 
valid during a READ, and done updating location during a WRITE */

// structural nets
wire [cam_depth_max-1:0] mbits0, mbits1, grp;
wire [md_max-1:0] MEMint_out, CACHE_out, CACHE_in; // 14-bit wide data signals for MM and cache 

// wire c0, c1, c2;                                   // clock signals generated by the PLL
wire mem_clk, cache_clk;

wire [cam_arg_max-3:0] dout0, dout1; // should be same as TAG bits used (using only 7-bits of TAG for now)
wire [ma_max-3:0] MEMint_address; // internal memory address port (using 12-bits for now instead of 14-bits)	

// registered nets
reg	[ma_max-3:0] MEMint_RDaddress, MEMint_WRaddress; // internal memory (using only 12-bits for now)

reg	we0, we1, WRint, writeback;	// address sources
reg	miss, wren, hit0, hit1; // hit0 and hit1 are used for debugging only

reg [cam_depth_max-1:0] replace = {cam_depth_max{1'b0}}; // for each location in CAM 

reg	[ca_max-1:0] CACHE_address; // cache memory address width {replace-bit, group-bits,word address bits} = 1+2+3=6

reg	[cam_arg_max-3:0] din0, din1; // should be same as TAG bits used (using only 7-bits of TAG for now)

reg	[t_cnt_max:0] transfer_count;

reg	[cam_depth_max-1:0] cam0_init, cam1_init; // Valid flag: to mark the first upload of a block of data to each cache block location

reg	[cam_depth_max-1:0] cam0_dirty_bit, cam1_dirty_bit; // to record if the block was ever written while in the cache

// grp_addrs_field is used to capture the value of the group address field
integer	grp_addrs_field;

// The PLL unit/block generates three clock phases to sequence all events
// dxp_pll_3_v	my_pll 	(Clock, c0, c1, c2);

// instantiate the CAM memories
av_CAM_v my_cam0 (
                  we0,
                  1'b1, 
                  din0, 
				  MEM_address[ma_max-3:5], //tag bits (using 7-bits instead of total of 9-bits )
				  MEM_address[4:3], // address bits for group
				  dout0,
				  mbits0         // match bits (1-bit for each location)
				  );
				  
av_CAM_v my_cam1 (
                  we1,
                  1'b1, 
                  din1, 
				  MEM_address[ma_max-3:5], 
				  MEM_address[4:3], 
				  dout1,
				  mbits1
				  );

// Main Memory RAM
assign mem_clk = WRint ? c2 : c1;  // READ access this is driven by the c1 phase of the clock, while for a WRITE access by c2.

assign MEMint_address = writeback ? MEMint_WRaddress : MEMint_RDaddress;

avRISC621_slave0_ram1 my_ram_slave0 (
                       MEMint_address[ma_max-3:0], // we are only using 12-bits for simulation purpose
                       ~mem_clk, 
					   CACHE_out, // data_in
					   WRint, 
					   MEMint_out  // data_out connected to CACHE_in (if hit and write)
					   );

// Cache memory as RAM	
assign cache_clk = WRint ? c1 : c2;	// opposite clocks wrt MM Write on c1 and Read on c2 

assign CACHE_in = ((hit0 || hit1) && WR) ? MEM_in : MEMint_out;

av_cache_v my_cache (
                     CACHE_address, // cache address width {replace-bit, group-bits,word address bits} = 1+2+3=6
					 ~cache_clk, 
					 CACHE_in, // data_in (14-bits)
					 wren, 
					 CACHE_out // data_out (14-bits)
					 );

assign MEM_out =  CACHE_out;

// This 2to4 decoder identifies the group being accessed
av_2to4_dec	my_dec	(MEM_address[4:3], grp);


//-------------------------------------------------------------------------------------------------------------------------------//

//------------------------------------------------CODE STARTS HERE--------------------------------------------------------------//

// memory subsystem "Control Unit"
/* MEM_address (memory address) = TAG=7-bit [11:5]| Group=2-bit [4:3]| Word=3-bit [2:0] */

wire c0_not;
assign c0_not = ~c0; // memory works at falling edge of processor clock i.e. rising edge of c0_not

always@(posedge c0_not)
begin
  if(Resetn == 0)
  begin
  miss = 1'b1;
  transfer_count = {(t_cnt_max + 1){1'b0}};
  replace = 4'b0000;
  we0 = 0;
  we1 = 0;
  hit0 = 0;
  hit1 = 0;
  Done = 0;
  WRint = 0;
  
  cam0_init[cam_depth_max-1:0] = {cam_depth_max{1'b0}};
  cam1_init[cam_depth_max-1:0] = {cam_depth_max{1'b0}};
  
  cam0_dirty_bit[cam_depth_max-1:0] = {cam_depth_max{1'b0}};
  cam1_dirty_bit[cam_depth_max-1:0] = {cam_depth_max{1'b0}};
  end

  else
  begin
    grp_addrs_field = MEM_address[4:3];
	
//----------------------------------------------------HIT condition-------------------------------------------------------------//
	if(miss == 0)
	begin
	  we0 = 0;
	  we1 = 0;
	  hit0 = 0;
	  hit1 = 0;
	  Done = 0;
	  WRint = 0;
	  wren = 0;
	  if(|(mbits0 & grp & cam0_init))
	  begin
	    CACHE_address = {1'b0, MEM_address[4:0]}; // [Group-bits,Word-bits], 1'b0 is track of replace
		if(WR == 1) // 2-w cache write
		begin
		  cam0_dirty_bit[grp_addrs_field] = 1;
		  wren = 1; // cache write 
		end 
		else begin
		  wren = 0;  // cache read
		end 
		hit0 = 1;
		Done = 1;
		replace[grp_addrs_field] = 1;
	  end 
	  else if(|(mbits1 & grp & cam1_init))
	  begin
	    CACHE_address = {1'b1, MEM_address[4:0]}; // why 1'b1??
		if(WR == 1)
		begin
		  cam1_dirty_bit[grp_addrs_field] = 1;
		  wren = 1;
		end 
		else begin
		  wren = 0;
		end 
		hit1 = 1;
		Done = 1;
		replace[grp_addrs_field] = 1'b0;
	  end
	  else begin
	    miss = 1'b1;
		transfer_count = {(t_cnt_max){1'b0}};
	  end 
	end 
	
//--------------------------WRITEBACK condition -- executed if dirty-bit for block to be replaced is set ------------------------//

	writeback = (miss &  
				((~replace[grp_addrs_field] & cam0_dirty_bit[grp_addrs_field]) 
				| (replace[grp_addrs_field] & cam1_dirty_bit[grp_addrs_field]))
				);
	if(writeback == 1)
	begin
	  wren = 0;
	  we0 = 0;
	  we1 = 0;
	  WRint = 1; // write to MM 
// replace[i] is 0 or 1, and is actually implementing a very simple replacement strategy: replace the 
// block that was not used last of the two blocks in the cache.
	  CACHE_address = {replace[grp_addrs_field], MEM_address[4:3], transfer_count[2:0]};
	  
	  if(replace[grp_addrs_field] == 0)
	    MEMint_WRaddress = {dout0, MEM_address[4:3], transfer_count[2:0]};
	  else
	    MEMint_WRaddress = {dout1, MEM_address[4:3], transfer_count[2:0]};
	  
	  transfer_count = transfer_count + 1'b1; // increment transfer count to point to next word in the block
	  if(transfer_count == 4'b1001)
	  begin
	    transfer_count = {(t_cnt_max+1){1'b0}}; // writeback = 1
		  if(replace[grp_addrs_field] == 0)
		    cam0_dirty_bit[grp_addrs_field] = 0;
		  else 
		    cam1_dirty_bit[grp_addrs_field] = 0;
	  end 
	end 
	
//------------------------------MISS condition -- upload requested block in the cache-----------------------------------------//

	if(miss == 1 && writeback == 0) begin
	CACHE_address = { replace[grp_addrs_field], MEM_address[4:3], transfer_count[2:0] };
	
	MEMint_RDaddress = {MEM_address[ma_max-3:3], transfer_count[2:0]};  // entire address generated by CPU 
	
	wren = 1; WRint = 0; // wren enables writing of next word into the cache 
	transfer_count = transfer_count + 1'b1; // increment the word transfer count to point to next word 
	
	if(transfer_count == 4'b1001)
	begin
	  miss = 0;
	  wren = 0;
	  transfer_count = 4'h0;
	  if(replace[grp_addrs_field] == 0)
	  begin
	    din0 = MEM_address[ma_max-3:5]; // TAG
		we0 = 1;
		if(cam0_init[grp_addrs_field] == 0)
		  cam0_init[grp_addrs_field] = 1;
	  end 
	  else begin
	    din1 = MEM_address[ma_max-3:5]; // TAG 
		we1 = 1;
		if(cam1_init[grp_addrs_field] == 0)
		  cam1_init[grp_addrs_field] = 1;
	  end 
	end 
	end
  
  end

end

endmodule



		  